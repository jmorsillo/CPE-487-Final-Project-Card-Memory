(paste code here)
