(Enter vga_sync.vhd)
