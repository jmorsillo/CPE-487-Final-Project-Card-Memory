(Put code here)
